-- megafunction wizard: %ALTPLL%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altpll 

-- ============================================================
-- File Name: vga_pll.vhd
-- Megafunction Name(s):
-- 			altpll
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 10.0 Build 262 08/18/2010 SP 1 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2010 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

Library UNISIM;
use UNISIM.vcomponents.all;

ENTITY vga_pll IS
	PORT
	(
		inclk0		: IN STD_LOGIC  := '0';
		c0		: OUT STD_LOGIC ;
		c1		: OUT STD_LOGIC 
	);
END vga_pll;

ARCHITECTURE SYN OF vga_pll IS
   signal clkfb : std_logic;
   signal clk25 : std_logic;
BEGIN
   c0 <= clkfb;
   c1 <= clk25;
   
   DCM_SP_inst : DCM_SP
   generic map (
      CLKDV_DIVIDE => 2.0,
      CLKFX_DIVIDE => 1,
      CLKFX_MULTIPLY => 2,
      CLKIN_DIVIDE_BY_2 => FALSE,
      CLKIN_PERIOD => 20.0, 
      CLKOUT_PHASE_SHIFT => "NONE", 
      CLK_FEEDBACK => "1X",         
      DESKEW_ADJUST => "SYSTEM_SYNCHRONOUS", 
      DLL_FREQUENCY_MODE => "LOW",
      DUTY_CYCLE_CORRECTION => TRUE, 
      PHASE_SHIFT => 0,        
      STARTUP_WAIT => FALSE) 
   port map (
      CLK0     => clkfb,     
      CLK180   => open, 
      CLK270   => open, -- 270 degree DCM CLK output
      CLK2X    => open,   -- 2X DCM CLK output
      CLK2X180 => open, -- 2X, 180 degree DCM CLK out
      CLK90    => open,   -- 90 degree DCM CLK output
      CLKDV    => clk25,   -- Divided DCM CLK out (CLKDV_DIVIDE)
      CLKFX    => open,   -- DCM CLK synthesis out (M/D)
      CLKFX180 => open, -- 180 degree CLK synthesis out
      LOCKED   => open, -- DCM LOCK status output
      PSDONE   => open, -- Dynamic phase adjust done output
      STATUS   => open, -- 8-bit DCM status bits output
      CLKFB    => CLKFB,   -- DCM clock feedback
      CLKIN    => inclk0,   -- Clock input (from IBUFG, BUFG or DCM)
      PSCLK    => '0',   -- Dynamic phase adjust clock input
      PSEN     => '0',     -- Dynamic phase adjust enable input
      PSINCDEC => '0', -- Dynamic phase adjust increment/decrement
      RST      => '0'        -- DCM asynchronous reset input
   );


END SYN;
